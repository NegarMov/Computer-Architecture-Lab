----------------------------------------------------------------------------------
-- Company:  		 AUT
-- Author: 			 Negar Movaghatian
-- Student ID:		 9831062
-- 
-- Create Date:    16:43:41 10/08/2021 
-- Design Name:    XOR Gate with 2 Inputs
-- Module Name:    xor_gate - Behavioral 
-- Project Name:   Computer Architecture Workshop 01
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity xor_gate is
    Port ( a : in  STD_LOGIC;
           b : in  STD_LOGIC;
           c : out  STD_LOGIC);
end xor_gate;

architecture Behavioral of xor_gate is

begin
	c <= a xor b;
	
end Behavioral;
